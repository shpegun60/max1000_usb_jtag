/******************* Power UP Reset Logic *********************/

module reset #(
	parameter logic RESET_OFF = 1'b1,                              // Defining a value of RESET
	parameter logic [24:0] POWER_UP_COUNTER_DELAY = 25'd25_000_000 // generate a 500ms reset pulse on initial powerup
)
(
  input  i_clk,
  output o_reset,
  output heart_bit
);

logic [24:0] PowUp_count = '0;        // counter reset
logic        PowUp_reset = ~RESET_OFF; // reset generated by
logic        toggle      = 1'b0;      // only for testing

// init values
initial begin
	PowUp_reset <= ~RESET_OFF; // reset generated by value
	toggle      <= 1'b0;
	PowUp_count <= '0;
end

always_ff @(posedge i_clk) begin
	PowUp_count <= PowUp_count + 1'b1;
	
	if (PowUp_count == POWER_UP_COUNTER_DELAY) begin 
		PowUp_reset <= RESET_OFF; 
		toggle      <= ~toggle;  // only for testing
	end
end

assign o_reset = PowUp_reset;

assign heart_bit = toggle;

endmodule
